`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:23:00 12/05/2018 
// Design Name: 
// Module Name:    mem_sin 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mem_sin(
    input wire clk, //系统时钟50MHz
    input wire memclk, //更新时钟
    input wire [1:0] memmode, //模式
    output reg [7:0] pout //定时输出锯齿波数字量
    );

// reg [19:0]cntdiv=0; //计数器，用于控制锯齿波数字量的变换时间
reg [7:0] addr = 0; //锯齿波数字量的地址，宽度为3
// wire [7:0] pout_wire;

// always@(posedge memclk) //计数器控制数字量输出的时间间隔
//     // if(cntdiv=='b101111101011110000) // 1Hz
//     if(cntdiv=='b11000011) //992Hz
//     begin
//         addr<=addr+1;
//         cntdiv<=1'b0;
//     end
//     else
//         cntdiv<=cntdiv+1'b1;

always@(posedge memclk) addr <= addr+1;

// rom_sin rom_sin(clk, addr, pout);

always@(posedge clk) //根据地址输出数字量
    if(memmode==2'b00) begin // Line
        pout<=8'b10000000;
        end
    else if(memmode==2'b01) begin // Triangular Wave
        pout <= addr;
        end
    else if(memmode==2'b10) begin // Square Wave
        case(addr[7])
            'b0:pout<=8'b11111111;
            'b1:pout<=8'b00000000;
        endcase
        end
    else if(memmode==2'b11) begin // Sine Wave
    case(addr)
        8'b00000000:pout<=8'b10000000;
        8'b00000001:pout<=8'b10000011;
        8'b00000010:pout<=8'b10000110;
        8'b00000011:pout<=8'b10001001;
        8'b00000100:pout<=8'b10001100;
        8'b00000101:pout<=8'b10001111;
        8'b00000110:pout<=8'b10010010;
        8'b00000111:pout<=8'b10010101;
        8'b00001000:pout<=8'b10011000;
        8'b00001001:pout<=8'b10011100;
        8'b00001010:pout<=8'b10011111;
        8'b00001011:pout<=8'b10100010;
        8'b00001100:pout<=8'b10100101;
        8'b00001101:pout<=8'b10101000;
        8'b00001110:pout<=8'b10101011;
        8'b00001111:pout<=8'b10101110;
        8'b00010000:pout<=8'b10110000;
        8'b00010001:pout<=8'b10110011;
        8'b00010010:pout<=8'b10110110;
        8'b00010011:pout<=8'b10111001;
        8'b00010100:pout<=8'b10111100;
        8'b00010101:pout<=8'b10111111;
        8'b00010110:pout<=8'b11000001;
        8'b00010111:pout<=8'b11000100;
        8'b00011000:pout<=8'b11000111;
        8'b00011001:pout<=8'b11001001;
        8'b00011010:pout<=8'b11001100;
        8'b00011011:pout<=8'b11001110;
        8'b00011100:pout<=8'b11010001;
        8'b00011101:pout<=8'b11010011;
        8'b00011110:pout<=8'b11010101;
        8'b00011111:pout<=8'b11011000;
        8'b00100000:pout<=8'b11011010;
        8'b00100001:pout<=8'b11011100;
        8'b00100010:pout<=8'b11011110;
        8'b00100011:pout<=8'b11100000;
        8'b00100100:pout<=8'b11100010;
        8'b00100101:pout<=8'b11100100;
        8'b00100110:pout<=8'b11100110;
        8'b00100111:pout<=8'b11101000;
        8'b00101000:pout<=8'b11101010;
        8'b00101001:pout<=8'b11101100;
        8'b00101010:pout<=8'b11101101;
        8'b00101011:pout<=8'b11101111;
        8'b00101100:pout<=8'b11110000;
        8'b00101101:pout<=8'b11110010;
        8'b00101110:pout<=8'b11110011;
        8'b00101111:pout<=8'b11110101;
        8'b00110000:pout<=8'b11110110;
        8'b00110001:pout<=8'b11110111;
        8'b00110010:pout<=8'b11111000;
        8'b00110011:pout<=8'b11111001;
        8'b00110100:pout<=8'b11111010;
        8'b00110101:pout<=8'b11111011;
        8'b00110110:pout<=8'b11111100;
        8'b00110111:pout<=8'b11111100;
        8'b00111000:pout<=8'b11111101;
        8'b00111001:pout<=8'b11111110;
        8'b00111010:pout<=8'b11111110;
        8'b00111011:pout<=8'b11111111;
        8'b00111100:pout<=8'b11111111;
        8'b00111101:pout<=8'b11111111;
        8'b00111110:pout<=8'b11111111;
        8'b00111111:pout<=8'b11111111;
        8'b01000000:pout<=8'b11111111;
        8'b01000001:pout<=8'b11111111;
        8'b01000010:pout<=8'b11111111;
        8'b01000011:pout<=8'b11111111;
        8'b01000100:pout<=8'b11111111;
        8'b01000101:pout<=8'b11111111;
        8'b01000110:pout<=8'b11111110;
        8'b01000111:pout<=8'b11111110;
        8'b01001000:pout<=8'b11111101;
        8'b01001001:pout<=8'b11111100;
        8'b01001010:pout<=8'b11111100;
        8'b01001011:pout<=8'b11111011;
        8'b01001100:pout<=8'b11111010;
        8'b01001101:pout<=8'b11111001;
        8'b01001110:pout<=8'b11111000;
        8'b01001111:pout<=8'b11110111;
        8'b01010000:pout<=8'b11110110;
        8'b01010001:pout<=8'b11110101;
        8'b01010010:pout<=8'b11110011;
        8'b01010011:pout<=8'b11110010;
        8'b01010100:pout<=8'b11110000;
        8'b01010101:pout<=8'b11101111;
        8'b01010110:pout<=8'b11101101;
        8'b01010111:pout<=8'b11101100;
        8'b01011000:pout<=8'b11101010;
        8'b01011001:pout<=8'b11101000;
        8'b01011010:pout<=8'b11100110;
        8'b01011011:pout<=8'b11100100;
        8'b01011100:pout<=8'b11100010;
        8'b01011101:pout<=8'b11100000;
        8'b01011110:pout<=8'b11011110;
        8'b01011111:pout<=8'b11011100;
        8'b01100000:pout<=8'b11011010;
        8'b01100001:pout<=8'b11011000;
        8'b01100010:pout<=8'b11010101;
        8'b01100011:pout<=8'b11010011;
        8'b01100100:pout<=8'b11010001;
        8'b01100101:pout<=8'b11001110;
        8'b01100110:pout<=8'b11001100;
        8'b01100111:pout<=8'b11001001;
        8'b01101000:pout<=8'b11000111;
        8'b01101001:pout<=8'b11000100;
        8'b01101010:pout<=8'b11000001;
        8'b01101011:pout<=8'b10111111;
        8'b01101100:pout<=8'b10111100;
        8'b01101101:pout<=8'b10111001;
        8'b01101110:pout<=8'b10110110;
        8'b01101111:pout<=8'b10110011;
        8'b01110000:pout<=8'b10110000;
        8'b01110001:pout<=8'b10101110;
        8'b01110010:pout<=8'b10101011;
        8'b01110011:pout<=8'b10101000;
        8'b01110100:pout<=8'b10100101;
        8'b01110101:pout<=8'b10100010;
        8'b01110110:pout<=8'b10011111;
        8'b01110111:pout<=8'b10011100;
        8'b01111000:pout<=8'b10011000;
        8'b01111001:pout<=8'b10010101;
        8'b01111010:pout<=8'b10010010;
        8'b01111011:pout<=8'b10001111;
        8'b01111100:pout<=8'b10001100;
        8'b01111101:pout<=8'b10001001;
        8'b01111110:pout<=8'b10000110;
        8'b01111111:pout<=8'b10000011;
        8'b10000000:pout<=8'b10000000;
        8'b10000001:pout<=8'b01111100;
        8'b10000010:pout<=8'b01111001;
        8'b10000011:pout<=8'b01110110;
        8'b10000100:pout<=8'b01110011;
        8'b10000101:pout<=8'b01110000;
        8'b10000110:pout<=8'b01101101;
        8'b10000111:pout<=8'b01101010;
        8'b10001000:pout<=8'b01100111;
        8'b10001001:pout<=8'b01100011;
        8'b10001010:pout<=8'b01100000;
        8'b10001011:pout<=8'b01011101;
        8'b10001100:pout<=8'b01011010;
        8'b10001101:pout<=8'b01010111;
        8'b10001110:pout<=8'b01010100;
        8'b10001111:pout<=8'b01010001;
        8'b10010000:pout<=8'b01001111;
        8'b10010001:pout<=8'b01001100;
        8'b10010010:pout<=8'b01001001;
        8'b10010011:pout<=8'b01000110;
        8'b10010100:pout<=8'b01000011;
        8'b10010101:pout<=8'b01000000;
        8'b10010110:pout<=8'b00111110;
        8'b10010111:pout<=8'b00111011;
        8'b10011000:pout<=8'b00111000;
        8'b10011001:pout<=8'b00110110;
        8'b10011010:pout<=8'b00110011;
        8'b10011011:pout<=8'b00110001;
        8'b10011100:pout<=8'b00101110;
        8'b10011101:pout<=8'b00101100;
        8'b10011110:pout<=8'b00101010;
        8'b10011111:pout<=8'b00100111;
        8'b10100000:pout<=8'b00100101;
        8'b10100001:pout<=8'b00100011;
        8'b10100010:pout<=8'b00100001;
        8'b10100011:pout<=8'b00011111;
        8'b10100100:pout<=8'b00011101;
        8'b10100101:pout<=8'b00011011;
        8'b10100110:pout<=8'b00011001;
        8'b10100111:pout<=8'b00010111;
        8'b10101000:pout<=8'b00010101;
        8'b10101001:pout<=8'b00010011;
        8'b10101010:pout<=8'b00010010;
        8'b10101011:pout<=8'b00010000;
        8'b10101100:pout<=8'b00001111;
        8'b10101101:pout<=8'b00001101;
        8'b10101110:pout<=8'b00001100;
        8'b10101111:pout<=8'b00001010;
        8'b10110000:pout<=8'b00001001;
        8'b10110001:pout<=8'b00001000;
        8'b10110010:pout<=8'b00000111;
        8'b10110011:pout<=8'b00000110;
        8'b10110100:pout<=8'b00000101;
        8'b10110101:pout<=8'b00000100;
        8'b10110110:pout<=8'b00000011;
        8'b10110111:pout<=8'b00000011;
        8'b10111000:pout<=8'b00000010;
        8'b10111001:pout<=8'b00000001;
        8'b10111010:pout<=8'b00000001;
        8'b10111011:pout<=8'b00000000;
        8'b10111100:pout<=8'b00000000;
        8'b10111101:pout<=8'b00000000;
        8'b10111110:pout<=8'b00000000;
        8'b10111111:pout<=8'b00000000;
        8'b11000000:pout<=8'b00000000;
        8'b11000001:pout<=8'b00000000;
        8'b11000010:pout<=8'b00000000;
        8'b11000011:pout<=8'b00000000;
        8'b11000100:pout<=8'b00000000;
        8'b11000101:pout<=8'b00000000;
        8'b11000110:pout<=8'b00000001;
        8'b11000111:pout<=8'b00000001;
        8'b11001000:pout<=8'b00000010;
        8'b11001001:pout<=8'b00000011;
        8'b11001010:pout<=8'b00000011;
        8'b11001011:pout<=8'b00000100;
        8'b11001100:pout<=8'b00000101;
        8'b11001101:pout<=8'b00000110;
        8'b11001110:pout<=8'b00000111;
        8'b11001111:pout<=8'b00001000;
        8'b11010000:pout<=8'b00001001;
        8'b11010001:pout<=8'b00001010;
        8'b11010010:pout<=8'b00001100;
        8'b11010011:pout<=8'b00001101;
        8'b11010100:pout<=8'b00001111;
        8'b11010101:pout<=8'b00010000;
        8'b11010110:pout<=8'b00010010;
        8'b11010111:pout<=8'b00010011;
        8'b11011000:pout<=8'b00010101;
        8'b11011001:pout<=8'b00010111;
        8'b11011010:pout<=8'b00011001;
        8'b11011011:pout<=8'b00011011;
        8'b11011100:pout<=8'b00011101;
        8'b11011101:pout<=8'b00011111;
        8'b11011110:pout<=8'b00100001;
        8'b11011111:pout<=8'b00100011;
        8'b11100000:pout<=8'b00100101;
        8'b11100001:pout<=8'b00100111;
        8'b11100010:pout<=8'b00101010;
        8'b11100011:pout<=8'b00101100;
        8'b11100100:pout<=8'b00101110;
        8'b11100101:pout<=8'b00110001;
        8'b11100110:pout<=8'b00110011;
        8'b11100111:pout<=8'b00110110;
        8'b11101000:pout<=8'b00111000;
        8'b11101001:pout<=8'b00111011;
        8'b11101010:pout<=8'b00111110;
        8'b11101011:pout<=8'b01000000;
        8'b11101100:pout<=8'b01000011;
        8'b11101101:pout<=8'b01000110;
        8'b11101110:pout<=8'b01001001;
        8'b11101111:pout<=8'b01001100;
        8'b11110000:pout<=8'b01001111;
        8'b11110001:pout<=8'b01010001;
        8'b11110010:pout<=8'b01010100;
        8'b11110011:pout<=8'b01010111;
        8'b11110100:pout<=8'b01011010;
        8'b11110101:pout<=8'b01011101;
        8'b11110110:pout<=8'b01100000;
        8'b11110111:pout<=8'b01100011;
        8'b11111000:pout<=8'b01100111;
        8'b11111001:pout<=8'b01101010;
        8'b11111010:pout<=8'b01101101;
        8'b11111011:pout<=8'b01110000;
        8'b11111100:pout<=8'b01110011;
        8'b11111101:pout<=8'b01110110;
        8'b11111110:pout<=8'b01111001;
        8'b11111111:pout<=8'b01111100;
        endcase
        end
endmodule
